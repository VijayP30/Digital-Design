`include "lab2_3_tb.sv"