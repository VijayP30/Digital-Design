`include "lab2_2_tb_file.sv"