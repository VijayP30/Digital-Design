`include "lab2_part1_tb.sv"