`include "Top_Level.sv"
`include "alarm.sv"
`include "ct_mod_N.sv"
`include "lcd_int3.sv"